// processador.v

// Generated using ACDS version 13.1 162 at 2018.08.08.12:34:48

`timescale 1 ps / 1 ps
module processador (
		input  wire        clk_clk,             //       clk.clk
		input  wire        reset_reset_n,       //     reset.reset_n
		output wire [3:0]  ledout_export,       //    ledout.export
		input  wire        botaoout_export,     //  botaoout.export
		output wire        wren_wren,           //      wren.wren
		output wire        data_data,           //      data.data
		output wire [31:0] wraddress_wraddress  // wraddress.wraddress
	);

	wire  [31:0] nios2_qsys_0_custom_instruction_master_result;                                  // nios2_qsys_0_custom_instruction_master_translator:ci_slave_result -> nios2_qsys_0:E_ci_result
	wire   [4:0] nios2_qsys_0_custom_instruction_master_b;                                       // nios2_qsys_0:D_ci_b -> nios2_qsys_0_custom_instruction_master_translator:ci_slave_b
	wire   [4:0] nios2_qsys_0_custom_instruction_master_c;                                       // nios2_qsys_0:D_ci_c -> nios2_qsys_0_custom_instruction_master_translator:ci_slave_c
	wire   [4:0] nios2_qsys_0_custom_instruction_master_a;                                       // nios2_qsys_0:D_ci_a -> nios2_qsys_0_custom_instruction_master_translator:ci_slave_a
	wire   [7:0] nios2_qsys_0_custom_instruction_master_n;                                       // nios2_qsys_0:D_ci_n -> nios2_qsys_0_custom_instruction_master_translator:ci_slave_n
	wire         nios2_qsys_0_custom_instruction_master_writerc;                                 // nios2_qsys_0:D_ci_writerc -> nios2_qsys_0_custom_instruction_master_translator:ci_slave_writerc
	wire  [31:0] nios2_qsys_0_custom_instruction_master_dataa;                                   // nios2_qsys_0:E_ci_dataa -> nios2_qsys_0_custom_instruction_master_translator:ci_slave_dataa
	wire         nios2_qsys_0_custom_instruction_master_readra;                                  // nios2_qsys_0:D_ci_readra -> nios2_qsys_0_custom_instruction_master_translator:ci_slave_readra
	wire  [31:0] nios2_qsys_0_custom_instruction_master_datab;                                   // nios2_qsys_0:E_ci_datab -> nios2_qsys_0_custom_instruction_master_translator:ci_slave_datab
	wire         nios2_qsys_0_custom_instruction_master_readrb;                                  // nios2_qsys_0:D_ci_readrb -> nios2_qsys_0_custom_instruction_master_translator:ci_slave_readrb
	wire  [31:0] nios2_qsys_0_custom_instruction_master_translator_comb_ci_master_result;        // nios2_qsys_0_custom_instruction_master_comb_xconnect:ci_slave_result -> nios2_qsys_0_custom_instruction_master_translator:comb_ci_master_result
	wire   [4:0] nios2_qsys_0_custom_instruction_master_translator_comb_ci_master_b;             // nios2_qsys_0_custom_instruction_master_translator:comb_ci_master_b -> nios2_qsys_0_custom_instruction_master_comb_xconnect:ci_slave_b
	wire   [4:0] nios2_qsys_0_custom_instruction_master_translator_comb_ci_master_c;             // nios2_qsys_0_custom_instruction_master_translator:comb_ci_master_c -> nios2_qsys_0_custom_instruction_master_comb_xconnect:ci_slave_c
	wire  [31:0] nios2_qsys_0_custom_instruction_master_translator_comb_ci_master_dataa;         // nios2_qsys_0_custom_instruction_master_translator:comb_ci_master_dataa -> nios2_qsys_0_custom_instruction_master_comb_xconnect:ci_slave_dataa
	wire   [4:0] nios2_qsys_0_custom_instruction_master_translator_comb_ci_master_a;             // nios2_qsys_0_custom_instruction_master_translator:comb_ci_master_a -> nios2_qsys_0_custom_instruction_master_comb_xconnect:ci_slave_a
	wire         nios2_qsys_0_custom_instruction_master_translator_comb_ci_master_readra;        // nios2_qsys_0_custom_instruction_master_translator:comb_ci_master_readra -> nios2_qsys_0_custom_instruction_master_comb_xconnect:ci_slave_readra
	wire   [7:0] nios2_qsys_0_custom_instruction_master_translator_comb_ci_master_n;             // nios2_qsys_0_custom_instruction_master_translator:comb_ci_master_n -> nios2_qsys_0_custom_instruction_master_comb_xconnect:ci_slave_n
	wire         nios2_qsys_0_custom_instruction_master_translator_comb_ci_master_writerc;       // nios2_qsys_0_custom_instruction_master_translator:comb_ci_master_writerc -> nios2_qsys_0_custom_instruction_master_comb_xconnect:ci_slave_writerc
	wire  [31:0] nios2_qsys_0_custom_instruction_master_translator_comb_ci_master_datab;         // nios2_qsys_0_custom_instruction_master_translator:comb_ci_master_datab -> nios2_qsys_0_custom_instruction_master_comb_xconnect:ci_slave_datab
	wire  [31:0] nios2_qsys_0_custom_instruction_master_translator_comb_ci_master_ipending;      // nios2_qsys_0_custom_instruction_master_translator:comb_ci_master_ipending -> nios2_qsys_0_custom_instruction_master_comb_xconnect:ci_slave_ipending
	wire         nios2_qsys_0_custom_instruction_master_translator_comb_ci_master_readrb;        // nios2_qsys_0_custom_instruction_master_translator:comb_ci_master_readrb -> nios2_qsys_0_custom_instruction_master_comb_xconnect:ci_slave_readrb
	wire         nios2_qsys_0_custom_instruction_master_translator_comb_ci_master_estatus;       // nios2_qsys_0_custom_instruction_master_translator:comb_ci_master_estatus -> nios2_qsys_0_custom_instruction_master_comb_xconnect:ci_slave_estatus
	wire  [31:0] nios2_qsys_0_custom_instruction_master_comb_xconnect_ci_master0_result;         // nios2_qsys_0_custom_instruction_master_comb_slave_translator0:ci_slave_result -> nios2_qsys_0_custom_instruction_master_comb_xconnect:ci_master0_result
	wire   [4:0] nios2_qsys_0_custom_instruction_master_comb_xconnect_ci_master0_b;              // nios2_qsys_0_custom_instruction_master_comb_xconnect:ci_master0_b -> nios2_qsys_0_custom_instruction_master_comb_slave_translator0:ci_slave_b
	wire   [4:0] nios2_qsys_0_custom_instruction_master_comb_xconnect_ci_master0_c;              // nios2_qsys_0_custom_instruction_master_comb_xconnect:ci_master0_c -> nios2_qsys_0_custom_instruction_master_comb_slave_translator0:ci_slave_c
	wire  [31:0] nios2_qsys_0_custom_instruction_master_comb_xconnect_ci_master0_dataa;          // nios2_qsys_0_custom_instruction_master_comb_xconnect:ci_master0_dataa -> nios2_qsys_0_custom_instruction_master_comb_slave_translator0:ci_slave_dataa
	wire   [4:0] nios2_qsys_0_custom_instruction_master_comb_xconnect_ci_master0_a;              // nios2_qsys_0_custom_instruction_master_comb_xconnect:ci_master0_a -> nios2_qsys_0_custom_instruction_master_comb_slave_translator0:ci_slave_a
	wire         nios2_qsys_0_custom_instruction_master_comb_xconnect_ci_master0_readra;         // nios2_qsys_0_custom_instruction_master_comb_xconnect:ci_master0_readra -> nios2_qsys_0_custom_instruction_master_comb_slave_translator0:ci_slave_readra
	wire   [7:0] nios2_qsys_0_custom_instruction_master_comb_xconnect_ci_master0_n;              // nios2_qsys_0_custom_instruction_master_comb_xconnect:ci_master0_n -> nios2_qsys_0_custom_instruction_master_comb_slave_translator0:ci_slave_n
	wire         nios2_qsys_0_custom_instruction_master_comb_xconnect_ci_master0_writerc;        // nios2_qsys_0_custom_instruction_master_comb_xconnect:ci_master0_writerc -> nios2_qsys_0_custom_instruction_master_comb_slave_translator0:ci_slave_writerc
	wire  [31:0] nios2_qsys_0_custom_instruction_master_comb_xconnect_ci_master0_datab;          // nios2_qsys_0_custom_instruction_master_comb_xconnect:ci_master0_datab -> nios2_qsys_0_custom_instruction_master_comb_slave_translator0:ci_slave_datab
	wire  [31:0] nios2_qsys_0_custom_instruction_master_comb_xconnect_ci_master0_ipending;       // nios2_qsys_0_custom_instruction_master_comb_xconnect:ci_master0_ipending -> nios2_qsys_0_custom_instruction_master_comb_slave_translator0:ci_slave_ipending
	wire         nios2_qsys_0_custom_instruction_master_comb_xconnect_ci_master0_readrb;         // nios2_qsys_0_custom_instruction_master_comb_xconnect:ci_master0_readrb -> nios2_qsys_0_custom_instruction_master_comb_slave_translator0:ci_slave_readrb
	wire         nios2_qsys_0_custom_instruction_master_comb_xconnect_ci_master0_estatus;        // nios2_qsys_0_custom_instruction_master_comb_xconnect:ci_master0_estatus -> nios2_qsys_0_custom_instruction_master_comb_slave_translator0:ci_slave_estatus
	wire  [31:0] nios2_qsys_0_custom_instruction_master_comb_slave_translator0_ci_master_result; // memoria_vga_0:result -> nios2_qsys_0_custom_instruction_master_comb_slave_translator0:ci_master_result
	wire  [31:0] nios2_qsys_0_custom_instruction_master_comb_slave_translator0_ci_master_dataa;  // nios2_qsys_0_custom_instruction_master_comb_slave_translator0:ci_master_dataa -> memoria_vga_0:dataa
	wire  [31:0] nios2_qsys_0_custom_instruction_master_comb_slave_translator0_ci_master_datab;  // nios2_qsys_0_custom_instruction_master_comb_slave_translator0:ci_master_datab -> memoria_vga_0:datab
	wire         mm_interconnect_0_nios2_qsys_0_jtag_debug_module_waitrequest;                   // nios2_qsys_0:jtag_debug_module_waitrequest -> mm_interconnect_0:nios2_qsys_0_jtag_debug_module_waitrequest
	wire  [31:0] mm_interconnect_0_nios2_qsys_0_jtag_debug_module_writedata;                     // mm_interconnect_0:nios2_qsys_0_jtag_debug_module_writedata -> nios2_qsys_0:jtag_debug_module_writedata
	wire   [8:0] mm_interconnect_0_nios2_qsys_0_jtag_debug_module_address;                       // mm_interconnect_0:nios2_qsys_0_jtag_debug_module_address -> nios2_qsys_0:jtag_debug_module_address
	wire         mm_interconnect_0_nios2_qsys_0_jtag_debug_module_write;                         // mm_interconnect_0:nios2_qsys_0_jtag_debug_module_write -> nios2_qsys_0:jtag_debug_module_write
	wire         mm_interconnect_0_nios2_qsys_0_jtag_debug_module_read;                          // mm_interconnect_0:nios2_qsys_0_jtag_debug_module_read -> nios2_qsys_0:jtag_debug_module_read
	wire  [31:0] mm_interconnect_0_nios2_qsys_0_jtag_debug_module_readdata;                      // nios2_qsys_0:jtag_debug_module_readdata -> mm_interconnect_0:nios2_qsys_0_jtag_debug_module_readdata
	wire         mm_interconnect_0_nios2_qsys_0_jtag_debug_module_debugaccess;                   // mm_interconnect_0:nios2_qsys_0_jtag_debug_module_debugaccess -> nios2_qsys_0:jtag_debug_module_debugaccess
	wire   [3:0] mm_interconnect_0_nios2_qsys_0_jtag_debug_module_byteenable;                    // mm_interconnect_0:nios2_qsys_0_jtag_debug_module_byteenable -> nios2_qsys_0:jtag_debug_module_byteenable
	wire  [31:0] mm_interconnect_0_onchip_memory2_0_s1_writedata;                                // mm_interconnect_0:onchip_memory2_0_s1_writedata -> onchip_memory2_0:writedata
	wire   [9:0] mm_interconnect_0_onchip_memory2_0_s1_address;                                  // mm_interconnect_0:onchip_memory2_0_s1_address -> onchip_memory2_0:address
	wire         mm_interconnect_0_onchip_memory2_0_s1_chipselect;                               // mm_interconnect_0:onchip_memory2_0_s1_chipselect -> onchip_memory2_0:chipselect
	wire         mm_interconnect_0_onchip_memory2_0_s1_clken;                                    // mm_interconnect_0:onchip_memory2_0_s1_clken -> onchip_memory2_0:clken
	wire         mm_interconnect_0_onchip_memory2_0_s1_write;                                    // mm_interconnect_0:onchip_memory2_0_s1_write -> onchip_memory2_0:write
	wire  [31:0] mm_interconnect_0_onchip_memory2_0_s1_readdata;                                 // onchip_memory2_0:readdata -> mm_interconnect_0:onchip_memory2_0_s1_readdata
	wire   [3:0] mm_interconnect_0_onchip_memory2_0_s1_byteenable;                               // mm_interconnect_0:onchip_memory2_0_s1_byteenable -> onchip_memory2_0:byteenable
	wire   [1:0] mm_interconnect_0_botao_s1_address;                                             // mm_interconnect_0:botao_s1_address -> botao:address
	wire  [31:0] mm_interconnect_0_botao_s1_readdata;                                            // botao:readdata -> mm_interconnect_0:botao_s1_readdata
	wire         nios2_qsys_0_data_master_waitrequest;                                           // mm_interconnect_0:nios2_qsys_0_data_master_waitrequest -> nios2_qsys_0:d_waitrequest
	wire  [31:0] nios2_qsys_0_data_master_writedata;                                             // nios2_qsys_0:d_writedata -> mm_interconnect_0:nios2_qsys_0_data_master_writedata
	wire  [13:0] nios2_qsys_0_data_master_address;                                               // nios2_qsys_0:d_address -> mm_interconnect_0:nios2_qsys_0_data_master_address
	wire         nios2_qsys_0_data_master_write;                                                 // nios2_qsys_0:d_write -> mm_interconnect_0:nios2_qsys_0_data_master_write
	wire         nios2_qsys_0_data_master_read;                                                  // nios2_qsys_0:d_read -> mm_interconnect_0:nios2_qsys_0_data_master_read
	wire  [31:0] nios2_qsys_0_data_master_readdata;                                              // mm_interconnect_0:nios2_qsys_0_data_master_readdata -> nios2_qsys_0:d_readdata
	wire         nios2_qsys_0_data_master_debugaccess;                                           // nios2_qsys_0:jtag_debug_module_debugaccess_to_roms -> mm_interconnect_0:nios2_qsys_0_data_master_debugaccess
	wire   [3:0] nios2_qsys_0_data_master_byteenable;                                            // nios2_qsys_0:d_byteenable -> mm_interconnect_0:nios2_qsys_0_data_master_byteenable
	wire  [31:0] mm_interconnect_0_leds_s1_writedata;                                            // mm_interconnect_0:leds_s1_writedata -> leds:writedata
	wire   [1:0] mm_interconnect_0_leds_s1_address;                                              // mm_interconnect_0:leds_s1_address -> leds:address
	wire         mm_interconnect_0_leds_s1_chipselect;                                           // mm_interconnect_0:leds_s1_chipselect -> leds:chipselect
	wire         mm_interconnect_0_leds_s1_write;                                                // mm_interconnect_0:leds_s1_write -> leds:write_n
	wire  [31:0] mm_interconnect_0_leds_s1_readdata;                                             // leds:readdata -> mm_interconnect_0:leds_s1_readdata
	wire         nios2_qsys_0_instruction_master_waitrequest;                                    // mm_interconnect_0:nios2_qsys_0_instruction_master_waitrequest -> nios2_qsys_0:i_waitrequest
	wire  [13:0] nios2_qsys_0_instruction_master_address;                                        // nios2_qsys_0:i_address -> mm_interconnect_0:nios2_qsys_0_instruction_master_address
	wire         nios2_qsys_0_instruction_master_read;                                           // nios2_qsys_0:i_read -> mm_interconnect_0:nios2_qsys_0_instruction_master_read
	wire  [31:0] nios2_qsys_0_instruction_master_readdata;                                       // mm_interconnect_0:nios2_qsys_0_instruction_master_readdata -> nios2_qsys_0:i_readdata
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest;                    // jtag_uart_0:av_waitrequest -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_waitrequest
	wire  [31:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata;                      // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_writedata -> jtag_uart_0:av_writedata
	wire   [0:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address;                        // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_address -> jtag_uart_0:av_address
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect;                     // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_chipselect -> jtag_uart_0:av_chipselect
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write;                          // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_write -> jtag_uart_0:av_write_n
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read;                           // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_read -> jtag_uart_0:av_read_n
	wire  [31:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata;                       // jtag_uart_0:av_readdata -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_readdata
	wire         irq_mapper_receiver0_irq;                                                       // jtag_uart_0:av_irq -> irq_mapper:receiver0_irq
	wire  [31:0] nios2_qsys_0_d_irq_irq;                                                         // irq_mapper:sender_irq -> nios2_qsys_0:d_irq
	wire         rst_controller_reset_out_reset;                                                 // rst_controller:reset_out -> [botao:reset_n, irq_mapper:reset, leds:reset_n, memoria_vga_0:reset, mm_interconnect_0:nios2_qsys_0_reset_n_reset_bridge_in_reset_reset, nios2_qsys_0:reset_n, onchip_memory2_0:reset, rst_translator:in_reset]
	wire         rst_controller_reset_out_reset_req;                                             // rst_controller:reset_req -> [nios2_qsys_0:reset_req, onchip_memory2_0:reset_req, rst_translator:reset_req_in]
	wire         rst_controller_001_reset_out_reset;                                             // rst_controller_001:reset_out -> [jtag_uart_0:rst_n, mm_interconnect_0:jtag_uart_0_reset_reset_bridge_in_reset_reset]
	wire         nios2_qsys_0_jtag_debug_module_reset_reset;                                     // nios2_qsys_0:jtag_debug_module_resetrequest -> rst_controller_001:reset_in0

	processador_nios2_qsys_0 nios2_qsys_0 (
		.clk                                   (clk_clk),                                                      //                       clk.clk
		.reset_n                               (~rst_controller_reset_out_reset),                              //                   reset_n.reset_n
		.reset_req                             (rst_controller_reset_out_reset_req),                           //                          .reset_req
		.d_address                             (nios2_qsys_0_data_master_address),                             //               data_master.address
		.d_byteenable                          (nios2_qsys_0_data_master_byteenable),                          //                          .byteenable
		.d_read                                (nios2_qsys_0_data_master_read),                                //                          .read
		.d_readdata                            (nios2_qsys_0_data_master_readdata),                            //                          .readdata
		.d_waitrequest                         (nios2_qsys_0_data_master_waitrequest),                         //                          .waitrequest
		.d_write                               (nios2_qsys_0_data_master_write),                               //                          .write
		.d_writedata                           (nios2_qsys_0_data_master_writedata),                           //                          .writedata
		.jtag_debug_module_debugaccess_to_roms (nios2_qsys_0_data_master_debugaccess),                         //                          .debugaccess
		.i_address                             (nios2_qsys_0_instruction_master_address),                      //        instruction_master.address
		.i_read                                (nios2_qsys_0_instruction_master_read),                         //                          .read
		.i_readdata                            (nios2_qsys_0_instruction_master_readdata),                     //                          .readdata
		.i_waitrequest                         (nios2_qsys_0_instruction_master_waitrequest),                  //                          .waitrequest
		.d_irq                                 (nios2_qsys_0_d_irq_irq),                                       //                     d_irq.irq
		.jtag_debug_module_resetrequest        (nios2_qsys_0_jtag_debug_module_reset_reset),                   //   jtag_debug_module_reset.reset
		.jtag_debug_module_address             (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_address),     //         jtag_debug_module.address
		.jtag_debug_module_byteenable          (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_byteenable),  //                          .byteenable
		.jtag_debug_module_debugaccess         (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_debugaccess), //                          .debugaccess
		.jtag_debug_module_read                (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_read),        //                          .read
		.jtag_debug_module_readdata            (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_readdata),    //                          .readdata
		.jtag_debug_module_waitrequest         (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_waitrequest), //                          .waitrequest
		.jtag_debug_module_write               (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_write),       //                          .write
		.jtag_debug_module_writedata           (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_writedata),   //                          .writedata
		.E_ci_result                           (nios2_qsys_0_custom_instruction_master_result),                // custom_instruction_master.result
		.D_ci_a                                (nios2_qsys_0_custom_instruction_master_a),                     //                          .a
		.D_ci_b                                (nios2_qsys_0_custom_instruction_master_b),                     //                          .b
		.D_ci_c                                (nios2_qsys_0_custom_instruction_master_c),                     //                          .c
		.D_ci_n                                (nios2_qsys_0_custom_instruction_master_n),                     //                          .n
		.D_ci_readra                           (nios2_qsys_0_custom_instruction_master_readra),                //                          .readra
		.D_ci_readrb                           (nios2_qsys_0_custom_instruction_master_readrb),                //                          .readrb
		.D_ci_writerc                          (nios2_qsys_0_custom_instruction_master_writerc),               //                          .writerc
		.E_ci_dataa                            (nios2_qsys_0_custom_instruction_master_dataa),                 //                          .dataa
		.E_ci_datab                            (nios2_qsys_0_custom_instruction_master_datab),                 //                          .datab
		.E_ci_multi_clock                      (),                                                             //                          .clk
		.E_ci_multi_reset                      (),                                                             //                          .reset
		.E_ci_multi_reset_req                  ()                                                              //                          .reset_req
	);

	processador_onchip_memory2_0 onchip_memory2_0 (
		.clk        (clk_clk),                                          //   clk1.clk
		.address    (mm_interconnect_0_onchip_memory2_0_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_onchip_memory2_0_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_onchip_memory2_0_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_onchip_memory2_0_s1_write),      //       .write
		.readdata   (mm_interconnect_0_onchip_memory2_0_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_onchip_memory2_0_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_onchip_memory2_0_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),                   // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req)                //       .reset_req
	);

	processador_leds leds (
		.clk        (clk_clk),                              //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address    (mm_interconnect_0_leds_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_leds_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_leds_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_leds_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_leds_s1_readdata),   //                    .readdata
		.out_port   (ledout_export)                         // external_connection.export
	);

	processador_botao botao (
		.clk      (clk_clk),                             //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),     //               reset.reset_n
		.address  (mm_interconnect_0_botao_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_botao_s1_readdata), //                    .readdata
		.in_port  (botaoout_export)                      // external_connection.export
	);

	processador_jtag_uart_0 jtag_uart_0 (
		.clk            (clk_clk),                                                     //               clk.clk
		.rst_n          (~rst_controller_001_reset_out_reset),                         //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver0_irq)                                     //               irq.irq
	);

	MSF #(
		.idle  (0),
		.faz   (1),
		.feito (2)
	) memoria_vga_0 (
		.clk       (clk_clk),                                                                        //                         clock.clk
		.reset     (rst_controller_reset_out_reset),                                                 //                         reset.reset
		.dataa     (nios2_qsys_0_custom_instruction_master_comb_slave_translator0_ci_master_dataa),  // nios_custom_instruction_slave.dataa
		.datab     (nios2_qsys_0_custom_instruction_master_comb_slave_translator0_ci_master_datab),  //                              .datab
		.result    (nios2_qsys_0_custom_instruction_master_comb_slave_translator0_ci_master_result), //                              .result
		.clken     (),                                                                               //                              .clk_en
		.start     (),                                                                               //                              .start
		.done      (),                                                                               //                              .done
		.wren      (wren_wren),                                                                      //                   conduit_end.wren
		.data      (data_data),                                                                      //                 conduit_end_1.data
		.wraddress (wraddress_wraddress)                                                             //                 conduit_end_2.wraddress
	);

	altera_customins_master_translator #(
		.SHARED_COMB_AND_MULTI (1)
	) nios2_qsys_0_custom_instruction_master_translator (
		.ci_slave_dataa            (nios2_qsys_0_custom_instruction_master_dataa),                              //       ci_slave.dataa
		.ci_slave_datab            (nios2_qsys_0_custom_instruction_master_datab),                              //               .datab
		.ci_slave_result           (nios2_qsys_0_custom_instruction_master_result),                             //               .result
		.ci_slave_n                (nios2_qsys_0_custom_instruction_master_n),                                  //               .n
		.ci_slave_readra           (nios2_qsys_0_custom_instruction_master_readra),                             //               .readra
		.ci_slave_readrb           (nios2_qsys_0_custom_instruction_master_readrb),                             //               .readrb
		.ci_slave_writerc          (nios2_qsys_0_custom_instruction_master_writerc),                            //               .writerc
		.ci_slave_a                (nios2_qsys_0_custom_instruction_master_a),                                  //               .a
		.ci_slave_b                (nios2_qsys_0_custom_instruction_master_b),                                  //               .b
		.ci_slave_c                (nios2_qsys_0_custom_instruction_master_c),                                  //               .c
		.ci_slave_ipending         (),                                                                          //               .ipending
		.ci_slave_estatus          (),                                                                          //               .estatus
		.comb_ci_master_dataa      (nios2_qsys_0_custom_instruction_master_translator_comb_ci_master_dataa),    // comb_ci_master.dataa
		.comb_ci_master_datab      (nios2_qsys_0_custom_instruction_master_translator_comb_ci_master_datab),    //               .datab
		.comb_ci_master_result     (nios2_qsys_0_custom_instruction_master_translator_comb_ci_master_result),   //               .result
		.comb_ci_master_n          (nios2_qsys_0_custom_instruction_master_translator_comb_ci_master_n),        //               .n
		.comb_ci_master_readra     (nios2_qsys_0_custom_instruction_master_translator_comb_ci_master_readra),   //               .readra
		.comb_ci_master_readrb     (nios2_qsys_0_custom_instruction_master_translator_comb_ci_master_readrb),   //               .readrb
		.comb_ci_master_writerc    (nios2_qsys_0_custom_instruction_master_translator_comb_ci_master_writerc),  //               .writerc
		.comb_ci_master_a          (nios2_qsys_0_custom_instruction_master_translator_comb_ci_master_a),        //               .a
		.comb_ci_master_b          (nios2_qsys_0_custom_instruction_master_translator_comb_ci_master_b),        //               .b
		.comb_ci_master_c          (nios2_qsys_0_custom_instruction_master_translator_comb_ci_master_c),        //               .c
		.comb_ci_master_ipending   (nios2_qsys_0_custom_instruction_master_translator_comb_ci_master_ipending), //               .ipending
		.comb_ci_master_estatus    (nios2_qsys_0_custom_instruction_master_translator_comb_ci_master_estatus),  //               .estatus
		.ci_slave_multi_clk        (1'b0),                                                                      //    (terminated)
		.ci_slave_multi_reset      (1'b0),                                                                      //    (terminated)
		.ci_slave_multi_clken      (1'b0),                                                                      //    (terminated)
		.ci_slave_multi_reset_req  (1'b0),                                                                      //    (terminated)
		.ci_slave_multi_start      (1'b0),                                                                      //    (terminated)
		.ci_slave_multi_done       (),                                                                          //    (terminated)
		.ci_slave_multi_dataa      (32'b00000000000000000000000000000000),                                      //    (terminated)
		.ci_slave_multi_datab      (32'b00000000000000000000000000000000),                                      //    (terminated)
		.ci_slave_multi_result     (),                                                                          //    (terminated)
		.ci_slave_multi_n          (8'b00000000),                                                               //    (terminated)
		.ci_slave_multi_readra     (1'b0),                                                                      //    (terminated)
		.ci_slave_multi_readrb     (1'b0),                                                                      //    (terminated)
		.ci_slave_multi_writerc    (1'b0),                                                                      //    (terminated)
		.ci_slave_multi_a          (5'b00000),                                                                  //    (terminated)
		.ci_slave_multi_b          (5'b00000),                                                                  //    (terminated)
		.ci_slave_multi_c          (5'b00000),                                                                  //    (terminated)
		.multi_ci_master_clk       (),                                                                          //    (terminated)
		.multi_ci_master_reset     (),                                                                          //    (terminated)
		.multi_ci_master_clken     (),                                                                          //    (terminated)
		.multi_ci_master_reset_req (),                                                                          //    (terminated)
		.multi_ci_master_start     (),                                                                          //    (terminated)
		.multi_ci_master_done      (1'b0),                                                                      //    (terminated)
		.multi_ci_master_dataa     (),                                                                          //    (terminated)
		.multi_ci_master_datab     (),                                                                          //    (terminated)
		.multi_ci_master_result    (32'b00000000000000000000000000000000),                                      //    (terminated)
		.multi_ci_master_n         (),                                                                          //    (terminated)
		.multi_ci_master_readra    (),                                                                          //    (terminated)
		.multi_ci_master_readrb    (),                                                                          //    (terminated)
		.multi_ci_master_writerc   (),                                                                          //    (terminated)
		.multi_ci_master_a         (),                                                                          //    (terminated)
		.multi_ci_master_b         (),                                                                          //    (terminated)
		.multi_ci_master_c         ()                                                                           //    (terminated)
	);

	processador_nios2_qsys_0_custom_instruction_master_comb_xconnect nios2_qsys_0_custom_instruction_master_comb_xconnect (
		.ci_slave_dataa      (nios2_qsys_0_custom_instruction_master_translator_comb_ci_master_dataa),    //   ci_slave.dataa
		.ci_slave_datab      (nios2_qsys_0_custom_instruction_master_translator_comb_ci_master_datab),    //           .datab
		.ci_slave_result     (nios2_qsys_0_custom_instruction_master_translator_comb_ci_master_result),   //           .result
		.ci_slave_n          (nios2_qsys_0_custom_instruction_master_translator_comb_ci_master_n),        //           .n
		.ci_slave_readra     (nios2_qsys_0_custom_instruction_master_translator_comb_ci_master_readra),   //           .readra
		.ci_slave_readrb     (nios2_qsys_0_custom_instruction_master_translator_comb_ci_master_readrb),   //           .readrb
		.ci_slave_writerc    (nios2_qsys_0_custom_instruction_master_translator_comb_ci_master_writerc),  //           .writerc
		.ci_slave_a          (nios2_qsys_0_custom_instruction_master_translator_comb_ci_master_a),        //           .a
		.ci_slave_b          (nios2_qsys_0_custom_instruction_master_translator_comb_ci_master_b),        //           .b
		.ci_slave_c          (nios2_qsys_0_custom_instruction_master_translator_comb_ci_master_c),        //           .c
		.ci_slave_ipending   (nios2_qsys_0_custom_instruction_master_translator_comb_ci_master_ipending), //           .ipending
		.ci_slave_estatus    (nios2_qsys_0_custom_instruction_master_translator_comb_ci_master_estatus),  //           .estatus
		.ci_master0_dataa    (nios2_qsys_0_custom_instruction_master_comb_xconnect_ci_master0_dataa),     // ci_master0.dataa
		.ci_master0_datab    (nios2_qsys_0_custom_instruction_master_comb_xconnect_ci_master0_datab),     //           .datab
		.ci_master0_result   (nios2_qsys_0_custom_instruction_master_comb_xconnect_ci_master0_result),    //           .result
		.ci_master0_n        (nios2_qsys_0_custom_instruction_master_comb_xconnect_ci_master0_n),         //           .n
		.ci_master0_readra   (nios2_qsys_0_custom_instruction_master_comb_xconnect_ci_master0_readra),    //           .readra
		.ci_master0_readrb   (nios2_qsys_0_custom_instruction_master_comb_xconnect_ci_master0_readrb),    //           .readrb
		.ci_master0_writerc  (nios2_qsys_0_custom_instruction_master_comb_xconnect_ci_master0_writerc),   //           .writerc
		.ci_master0_a        (nios2_qsys_0_custom_instruction_master_comb_xconnect_ci_master0_a),         //           .a
		.ci_master0_b        (nios2_qsys_0_custom_instruction_master_comb_xconnect_ci_master0_b),         //           .b
		.ci_master0_c        (nios2_qsys_0_custom_instruction_master_comb_xconnect_ci_master0_c),         //           .c
		.ci_master0_ipending (nios2_qsys_0_custom_instruction_master_comb_xconnect_ci_master0_ipending),  //           .ipending
		.ci_master0_estatus  (nios2_qsys_0_custom_instruction_master_comb_xconnect_ci_master0_estatus)    //           .estatus
	);

	altera_customins_slave_translator #(
		.N_WIDTH          (8),
		.USE_DONE         (1),
		.NUM_FIXED_CYCLES (0)
	) nios2_qsys_0_custom_instruction_master_comb_slave_translator0 (
		.ci_slave_dataa      (nios2_qsys_0_custom_instruction_master_comb_xconnect_ci_master0_dataa),          //  ci_slave.dataa
		.ci_slave_datab      (nios2_qsys_0_custom_instruction_master_comb_xconnect_ci_master0_datab),          //          .datab
		.ci_slave_result     (nios2_qsys_0_custom_instruction_master_comb_xconnect_ci_master0_result),         //          .result
		.ci_slave_n          (nios2_qsys_0_custom_instruction_master_comb_xconnect_ci_master0_n),              //          .n
		.ci_slave_readra     (nios2_qsys_0_custom_instruction_master_comb_xconnect_ci_master0_readra),         //          .readra
		.ci_slave_readrb     (nios2_qsys_0_custom_instruction_master_comb_xconnect_ci_master0_readrb),         //          .readrb
		.ci_slave_writerc    (nios2_qsys_0_custom_instruction_master_comb_xconnect_ci_master0_writerc),        //          .writerc
		.ci_slave_a          (nios2_qsys_0_custom_instruction_master_comb_xconnect_ci_master0_a),              //          .a
		.ci_slave_b          (nios2_qsys_0_custom_instruction_master_comb_xconnect_ci_master0_b),              //          .b
		.ci_slave_c          (nios2_qsys_0_custom_instruction_master_comb_xconnect_ci_master0_c),              //          .c
		.ci_slave_ipending   (nios2_qsys_0_custom_instruction_master_comb_xconnect_ci_master0_ipending),       //          .ipending
		.ci_slave_estatus    (nios2_qsys_0_custom_instruction_master_comb_xconnect_ci_master0_estatus),        //          .estatus
		.ci_master_dataa     (nios2_qsys_0_custom_instruction_master_comb_slave_translator0_ci_master_dataa),  // ci_master.dataa
		.ci_master_datab     (nios2_qsys_0_custom_instruction_master_comb_slave_translator0_ci_master_datab),  //          .datab
		.ci_master_result    (nios2_qsys_0_custom_instruction_master_comb_slave_translator0_ci_master_result), //          .result
		.ci_master_n         (),                                                                               // (terminated)
		.ci_master_readra    (),                                                                               // (terminated)
		.ci_master_readrb    (),                                                                               // (terminated)
		.ci_master_writerc   (),                                                                               // (terminated)
		.ci_master_a         (),                                                                               // (terminated)
		.ci_master_b         (),                                                                               // (terminated)
		.ci_master_c         (),                                                                               // (terminated)
		.ci_master_ipending  (),                                                                               // (terminated)
		.ci_master_estatus   (),                                                                               // (terminated)
		.ci_master_clk       (),                                                                               // (terminated)
		.ci_master_clken     (),                                                                               // (terminated)
		.ci_master_reset_req (),                                                                               // (terminated)
		.ci_master_reset     (),                                                                               // (terminated)
		.ci_master_start     (),                                                                               // (terminated)
		.ci_master_done      (1'b0),                                                                           // (terminated)
		.ci_slave_clk        (1'b0),                                                                           // (terminated)
		.ci_slave_clken      (1'b0),                                                                           // (terminated)
		.ci_slave_reset_req  (1'b0),                                                                           // (terminated)
		.ci_slave_reset      (1'b0),                                                                           // (terminated)
		.ci_slave_start      (1'b0),                                                                           // (terminated)
		.ci_slave_done       ()                                                                                // (terminated)
	);

	processador_mm_interconnect_0 mm_interconnect_0 (
		.clk_0_clk_clk                                    (clk_clk),                                                      //                                  clk_0_clk.clk
		.jtag_uart_0_reset_reset_bridge_in_reset_reset    (rst_controller_001_reset_out_reset),                           //    jtag_uart_0_reset_reset_bridge_in_reset.reset
		.nios2_qsys_0_reset_n_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                               // nios2_qsys_0_reset_n_reset_bridge_in_reset.reset
		.nios2_qsys_0_data_master_address                 (nios2_qsys_0_data_master_address),                             //                   nios2_qsys_0_data_master.address
		.nios2_qsys_0_data_master_waitrequest             (nios2_qsys_0_data_master_waitrequest),                         //                                           .waitrequest
		.nios2_qsys_0_data_master_byteenable              (nios2_qsys_0_data_master_byteenable),                          //                                           .byteenable
		.nios2_qsys_0_data_master_read                    (nios2_qsys_0_data_master_read),                                //                                           .read
		.nios2_qsys_0_data_master_readdata                (nios2_qsys_0_data_master_readdata),                            //                                           .readdata
		.nios2_qsys_0_data_master_write                   (nios2_qsys_0_data_master_write),                               //                                           .write
		.nios2_qsys_0_data_master_writedata               (nios2_qsys_0_data_master_writedata),                           //                                           .writedata
		.nios2_qsys_0_data_master_debugaccess             (nios2_qsys_0_data_master_debugaccess),                         //                                           .debugaccess
		.nios2_qsys_0_instruction_master_address          (nios2_qsys_0_instruction_master_address),                      //            nios2_qsys_0_instruction_master.address
		.nios2_qsys_0_instruction_master_waitrequest      (nios2_qsys_0_instruction_master_waitrequest),                  //                                           .waitrequest
		.nios2_qsys_0_instruction_master_read             (nios2_qsys_0_instruction_master_read),                         //                                           .read
		.nios2_qsys_0_instruction_master_readdata         (nios2_qsys_0_instruction_master_readdata),                     //                                           .readdata
		.botao_s1_address                                 (mm_interconnect_0_botao_s1_address),                           //                                   botao_s1.address
		.botao_s1_readdata                                (mm_interconnect_0_botao_s1_readdata),                          //                                           .readdata
		.jtag_uart_0_avalon_jtag_slave_address            (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address),      //              jtag_uart_0_avalon_jtag_slave.address
		.jtag_uart_0_avalon_jtag_slave_write              (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write),        //                                           .write
		.jtag_uart_0_avalon_jtag_slave_read               (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read),         //                                           .read
		.jtag_uart_0_avalon_jtag_slave_readdata           (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata),     //                                           .readdata
		.jtag_uart_0_avalon_jtag_slave_writedata          (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata),    //                                           .writedata
		.jtag_uart_0_avalon_jtag_slave_waitrequest        (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest),  //                                           .waitrequest
		.jtag_uart_0_avalon_jtag_slave_chipselect         (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect),   //                                           .chipselect
		.leds_s1_address                                  (mm_interconnect_0_leds_s1_address),                            //                                    leds_s1.address
		.leds_s1_write                                    (mm_interconnect_0_leds_s1_write),                              //                                           .write
		.leds_s1_readdata                                 (mm_interconnect_0_leds_s1_readdata),                           //                                           .readdata
		.leds_s1_writedata                                (mm_interconnect_0_leds_s1_writedata),                          //                                           .writedata
		.leds_s1_chipselect                               (mm_interconnect_0_leds_s1_chipselect),                         //                                           .chipselect
		.nios2_qsys_0_jtag_debug_module_address           (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_address),     //             nios2_qsys_0_jtag_debug_module.address
		.nios2_qsys_0_jtag_debug_module_write             (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_write),       //                                           .write
		.nios2_qsys_0_jtag_debug_module_read              (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_read),        //                                           .read
		.nios2_qsys_0_jtag_debug_module_readdata          (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_readdata),    //                                           .readdata
		.nios2_qsys_0_jtag_debug_module_writedata         (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_writedata),   //                                           .writedata
		.nios2_qsys_0_jtag_debug_module_byteenable        (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_byteenable),  //                                           .byteenable
		.nios2_qsys_0_jtag_debug_module_waitrequest       (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_waitrequest), //                                           .waitrequest
		.nios2_qsys_0_jtag_debug_module_debugaccess       (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_debugaccess), //                                           .debugaccess
		.onchip_memory2_0_s1_address                      (mm_interconnect_0_onchip_memory2_0_s1_address),                //                        onchip_memory2_0_s1.address
		.onchip_memory2_0_s1_write                        (mm_interconnect_0_onchip_memory2_0_s1_write),                  //                                           .write
		.onchip_memory2_0_s1_readdata                     (mm_interconnect_0_onchip_memory2_0_s1_readdata),               //                                           .readdata
		.onchip_memory2_0_s1_writedata                    (mm_interconnect_0_onchip_memory2_0_s1_writedata),              //                                           .writedata
		.onchip_memory2_0_s1_byteenable                   (mm_interconnect_0_onchip_memory2_0_s1_byteenable),             //                                           .byteenable
		.onchip_memory2_0_s1_chipselect                   (mm_interconnect_0_onchip_memory2_0_s1_chipselect),             //                                           .chipselect
		.onchip_memory2_0_s1_clken                        (mm_interconnect_0_onchip_memory2_0_s1_clken)                   //                                           .clken
	);

	processador_irq_mapper irq_mapper (
		.clk           (clk_clk),                        //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.sender_irq    (nios2_qsys_0_d_irq_irq)          //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (nios2_qsys_0_jtag_debug_module_reset_reset), // reset_in0.reset
		.reset_in1      (~reset_reset_n),                             // reset_in1.reset
		.clk            (clk_clk),                                    //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset),         // reset_out.reset
		.reset_req      (),                                           // (terminated)
		.reset_req_in0  (1'b0),                                       // (terminated)
		.reset_req_in1  (1'b0),                                       // (terminated)
		.reset_in2      (1'b0),                                       // (terminated)
		.reset_req_in2  (1'b0),                                       // (terminated)
		.reset_in3      (1'b0),                                       // (terminated)
		.reset_req_in3  (1'b0),                                       // (terminated)
		.reset_in4      (1'b0),                                       // (terminated)
		.reset_req_in4  (1'b0),                                       // (terminated)
		.reset_in5      (1'b0),                                       // (terminated)
		.reset_req_in5  (1'b0),                                       // (terminated)
		.reset_in6      (1'b0),                                       // (terminated)
		.reset_req_in6  (1'b0),                                       // (terminated)
		.reset_in7      (1'b0),                                       // (terminated)
		.reset_req_in7  (1'b0),                                       // (terminated)
		.reset_in8      (1'b0),                                       // (terminated)
		.reset_req_in8  (1'b0),                                       // (terminated)
		.reset_in9      (1'b0),                                       // (terminated)
		.reset_req_in9  (1'b0),                                       // (terminated)
		.reset_in10     (1'b0),                                       // (terminated)
		.reset_req_in10 (1'b0),                                       // (terminated)
		.reset_in11     (1'b0),                                       // (terminated)
		.reset_req_in11 (1'b0),                                       // (terminated)
		.reset_in12     (1'b0),                                       // (terminated)
		.reset_req_in12 (1'b0),                                       // (terminated)
		.reset_in13     (1'b0),                                       // (terminated)
		.reset_req_in13 (1'b0),                                       // (terminated)
		.reset_in14     (1'b0),                                       // (terminated)
		.reset_req_in14 (1'b0),                                       // (terminated)
		.reset_in15     (1'b0),                                       // (terminated)
		.reset_req_in15 (1'b0)                                        // (terminated)
	);

endmodule
