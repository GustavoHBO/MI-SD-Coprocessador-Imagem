// dma_controller.v

// Generated using ACDS version 13.1 162 at 2018.08.03.13:01:26

`timescale 1 ps / 1 ps
module dma_controller (
		input  wire        clk_clk,            //      clk.clk
		input  wire        reset_reset_n,      //    reset.reset_n
		input  wire [10:0] s2_port_address,    //  s2_port.address
		input  wire        s2_port_chipselect, //         .chipselect
		input  wire        s2_port_clken,      //         .clken
		input  wire        s2_port_write,      //         .write
		output wire [31:0] s2_port_readdata,   //         .readdata
		input  wire [31:0] s2_port_writedata,  //         .writedata
		input  wire [3:0]  s2_port_byteenable, //         .byteenable
		input  wire        s2_reset_reset,     // s2_reset.reset
		input  wire        s2_reset_reset_req  //         .reset_req
	);

	wire    rst_controller_reset_out_reset;     // rst_controller:reset_out -> onchip_memory2_0:reset
	wire    rst_controller_reset_out_reset_req; // rst_controller:reset_req -> onchip_memory2_0:reset_req

	dma_controller_onchip_memory2_0 onchip_memory2_0 (
		.clk         (clk_clk),                            //   clk1.clk
		.address     (),                                   //     s1.address
		.debugaccess (),                                   //       .debugaccess
		.clken       (),                                   //       .clken
		.chipselect  (),                                   //       .chipselect
		.write       (),                                   //       .write
		.readdata    (),                                   //       .readdata
		.writedata   (),                                   //       .writedata
		.byteenable  (),                                   //       .byteenable
		.reset       (rst_controller_reset_out_reset),     // reset1.reset
		.reset_req   (rst_controller_reset_out_reset_req), //       .reset_req
		.address2    (s2_port_address),                    //     s2.address
		.chipselect2 (s2_port_chipselect),                 //       .chipselect
		.clken2      (s2_port_clken),                      //       .clken
		.write2      (s2_port_write),                      //       .write
		.readdata2   (s2_port_readdata),                   //       .readdata
		.writedata2  (s2_port_writedata),                  //       .writedata
		.byteenable2 (s2_port_byteenable),                 //       .byteenable
		.clk2        (clk_clk),                            //   clk2.clk
		.reset2      (s2_reset_reset),                     // reset2.reset
		.reset_req2  (s2_reset_reset_req)                  //       .reset_req
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
