//------------------------------------------------------------------------------
//	Module:		Lab2Lock
//	Desc:			This module implements the functionality of a simple combination lock.
//					The lock uses 2 4-bit combination digits.
//					See the lab document for the suggested combination setting.
//	Params:		This module is not parameterized.
//	Inputs:		See Lab2 document
//	Outputs:	See Lab2 document
//
//	Author:     YOUR NAME GOES HERE
//------------------------------------------------------------------------------
module	Lab2Lock(
			//------------------------------------------------------------------
			//	Clock & Reset Inputs
			//------------------------------------------------------------------
			Clock,
			Reset,
			//------------------------------------------------------------------
			
			//------------------------------------------------------------------
			//	Inputs
			//------------------------------------------------------------------
			Enter,
			Digit,
			//------------------------------------------------------------------
			
			//------------------------------------------------------------------
			//	Outputs
			//------------------------------------------------------------------
			State,
			Open,
			Fail
			//------------------------------------------------------------------
	);
	//--------------------------------------------------------------------------
	//	Parameters
	//--------------------------------------------------------------------------
	localparam	DIGIT_1	=	4'h2,
					DIGIT_2	=	4'h3;
										
	//--------------------------------------------------------------------------
	
	//--------------------------------------------------------------------------
	//	Clock & Reset Inputs
	//--------------------------------------------------------------------------
	input					Clock;	// System clock
	input					Reset;	// System reset
	//--------------------------------------------------------------------------
	
	//--------------------------------------------------------------------------
	//	Inputs
	//--------------------------------------------------------------------------
	input					Enter;
	input		[3:0]		Digit;
	//--------------------------------------------------------------------------
	
	//--------------------------------------------------------------------------
	//	Outputs
	//--------------------------------------------------------------------------
	output	[2:0]		State;
	output	reg				Open;
	output	reg				Fail;
	//--------------------------------------------------------------------------

	//--------------------------------------------------------------------------
	//	State Encoding
	//--------------------------------------------------------------------------
	
	parameter [2:0] 	IDLE = 3'b000,
							LOCKED = 3'b001,
							BAD1 = 3'b011,
							BAD2 = 3'b010,
							OK = 3'b110,
							OPEN = 3'b111;
	
	// place state encoding here
	
	//--------------------------------------------------------------------------
	
	//--------------------------------------------------------------------------
	//	Wire Declarations
	//--------------------------------------------------------------------------
	
	// place wire declarations here	
	
	//--------------------------------------------------------------------------
	
	//--------------------------------------------------------------------------
	//	Logic
	//--------------------------------------------------------------------------
	
	// Place you *behavioral* Verilog here
	// You may find it useful to use a case statement to describe your FSM.
	
	reg [2:0] state, next;
	
	always @(posedge Clock) begin
		if (Reset) begin 
			state <= IDLE;
		end
		else begin 
			state <= next;
		end
	end
	assign State = state;
	
	always @(Enter or state) begin // Sempre que isso ocorrer, execute o codigo abaixo!
		case (state)
			IDLE : begin
				next = LOCKED;
				Open = 1'b0;
				Fail = 1'b0;
			end
			LOCKED : begin
				if(Enter) begin
					if (Digit == DIGIT_1) next = OK;
					else next = BAD1;
				end
				else next = LOCKED;
			end
			OK : begin
				if(Enter) begin
					if (Digit == DIGIT_2) next = OPEN;
					else next = BAD2;
				end
				else next = OK;
			end
			BAD1 : begin 
				if (Enter) next = BAD2;
				else next = BAD1;
			end
			BAD2 : begin 
				Fail = 1'b1;
				next = BAD2;
			end
			OPEN : begin 
				Open = 1'b1;
				next = OPEN;
			end
		endcase
	end
	
	//--------------------------------------------------------------------------
endmodule
//------------------------------------------------------------------------------
