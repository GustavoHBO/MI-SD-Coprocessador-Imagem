module convolution(
	input clk_in, 
	input [63:0]matrix_in,
	output [7:0]pixel_out
);

	output = 

endmodule 